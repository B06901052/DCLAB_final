timeunit		1ns;
timeprecision	1ns;

module GameController (
	input		i_clk,
	input		i_rst_n,
	input [1:0] i_mode,//0~2:1P easy, normal, hard; 3:2P
	input		i_start,
	input		i_surrender,
	input 		i_prestep,
);

/*================================================================*
 * LOCALPARAM
 *================================================================*/
localparam S_IDLE = 0;

/*================================================================*
 * REG/WIRE
 *================================================================*/
logic	state_r;

/*================================================================*
 * ASSIGN
 *================================================================*/

/*================================================================*
 * Sequential (state)
 *================================================================*/ 
always_ff @(posedge i_clk or negedge i_rst_n) begin
	if (!i_rst_n) begin
		state_r	<= S_IDLE;
	end else begin
		case (state_r)
		S_IDLE:begin
		
		end
		default:begin
		
		end
		endcase
	end
end

/*================================================================* 
 * Combination
 *================================================================*/ 
always_comb begin
	
end

/*================================================================* 
 * Module 
 *================================================================*/

endmodule